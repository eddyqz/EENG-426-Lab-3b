magic
tech sky130l
timestamp 1668056821
<< checkpaint >>
rect 48 40 113 105
<< error_s >>
rect 537 965 539 967
rect 596 964 598 966
rect 660 964 662 966
rect 745 965 747 967
rect 801 965 803 967
rect 376 899 378 902
rect 528 899 530 902
rect 648 899 650 902
rect 379 876 381 899
rect 531 876 533 899
rect 651 876 653 899
rect 664 827 668 828
rect 696 827 700 828
rect 760 827 764 828
rect 792 827 796 828
rect 504 807 506 810
rect 507 784 509 807
rect 722 789 725 790
rect 811 784 813 790
rect 717 770 722 771
rect 783 770 791 771
rect 754 649 757 650
rect 843 644 845 650
rect 744 636 748 637
rect 832 636 836 637
rect 741 630 751 631
rect 837 630 842 631
rect 432 620 434 623
rect 343 617 346 618
rect 435 617 437 620
rect 663 617 666 618
rect 250 537 253 538
rect 338 537 341 538
rect 247 449 250 450
rect 567 449 570 450
rect 655 449 658 450
rect 743 449 746 450
rect 831 449 834 450
rect 215 289 218 290
rect 303 289 306 290
rect 391 289 394 290
rect 479 289 482 290
rect 218 209 221 210
<< m2 >>
rect 300 1006 308 1008
rect 532 1006 540 1008
rect 756 1006 764 1008
rect 80 928 82 936
rect 982 920 984 928
rect 80 848 82 856
rect 982 832 984 840
rect 80 772 82 780
rect 982 748 984 756
rect 80 692 82 700
rect 982 664 984 672
rect 80 616 82 624
rect 982 580 984 588
rect 80 536 82 544
rect 982 492 984 500
rect 80 460 82 468
rect 982 408 984 416
rect 80 380 82 388
rect 982 324 984 332
rect 80 304 82 312
rect 982 240 984 248
rect 80 224 82 232
rect 80 148 82 156
rect 982 152 984 160
use circuitwell  npwells
timestamp 1668056821
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 1668056821
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1667968642
transform 1 0 104 0 1 92
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_alainv
timestamp 1668054752
transform 1 0 128 0 1 88
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_alainv
timestamp 1668054752
transform 1 0 160 0 1 88
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_alainv
timestamp 1668054752
transform 1 0 192 0 1 88
box 3 -1 28 37
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_55_6
timestamp 1667968642
transform 1 0 288 0 1 84
box 8 4 76 44
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_55_6
timestamp 1667968642
transform 1 0 256 0 1 88
box 8 4 28 36
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_55_6
timestamp 1668054752
transform 1 0 224 0 1 88
box 3 -1 28 37
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_55_6_anx
timestamp 1667968642
transform 1 0 368 0 1 84
box 8 4 36 60
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_55_6_al
timestamp 1667968642
transform 1 0 408 0 1 84
box 8 4 76 48
use _0_0std_0_0cells_0_0FAX1  add_afa_54_6
timestamp 1667968642
transform 1 0 488 0 1 76
box 8 4 140 84
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_54_6
timestamp 1667968642
transform 1 0 704 0 1 84
box 8 4 76 44
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_54_6_anx
timestamp 1667968642
transform 1 0 632 0 1 84
box 8 4 36 60
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_54_6
timestamp 1668054752
transform 1 0 672 0 1 88
box 3 -1 28 37
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_53_6
timestamp 1667968642
transform 1 0 856 0 1 84
box 8 4 76 44
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_53_6_anx
timestamp 1667968642
transform 1 0 816 0 1 84
box 8 4 36 60
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_53_6
timestamp 1668054752
transform 1 0 784 0 1 88
box 3 -1 28 37
use welltap_svt  __well_tap__1
timestamp 1667968642
transform 1 0 944 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1667968642
transform 1 0 104 0 -1 236
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_55_6
timestamp 1668056734
transform 1 0 128 0 -1 244
box 2 -1 90 54
use _0_0std_0_0cells_0_0FAX1  add_afa_55_6
timestamp 1667968642
transform 1 0 304 0 -1 252
box 8 4 140 84
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_54_6
timestamp 1668056734
transform 1 0 216 0 -1 244
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_54_6_al
timestamp 1667968642
transform 1 0 448 0 -1 244
box 8 4 76 48
use _0_0std_0_0cells_0_0FAX1  add_afa_53_6
timestamp 1667968642
transform 1 0 536 0 -1 252
box 8 4 140 84
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_54_6
timestamp 1667968642
transform 1 0 688 0 -1 240
box 8 4 28 36
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_53_6
timestamp 1668056734
transform 1 0 728 0 -1 244
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_53_6_al
timestamp 1667968642
transform 1 0 824 0 -1 244
box 8 4 76 48
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_53_6
timestamp 1667968642
transform 1 0 904 0 -1 240
box 8 4 28 36
use welltap_svt  __well_tap__3
timestamp 1667968642
transform 1 0 944 0 -1 236
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1667968642
transform 1 0 104 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_55_6
timestamp 1668056734
transform 1 0 128 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_55_6
timestamp 1668056734
transform 1 0 304 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_54_6
timestamp 1668056734
transform 1 0 216 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_54_6
timestamp 1668056734
transform 1 0 392 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_54_6
timestamp 1668056734
transform 1 0 480 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_53_6
timestamp 1668056734
transform 1 0 576 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_53_6
timestamp 1668056734
transform 1 0 672 0 1 252
box 2 -1 90 54
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_52_6_anx
timestamp 1667968642
transform 1 0 864 0 1 252
box 8 4 36 60
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_53_6
timestamp 1668056734
transform 1 0 768 0 1 252
box 2 -1 90 54
use welltap_svt  __well_tap__5
timestamp 1667968642
transform 1 0 944 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_57_6
timestamp 1667968642
transform 1 0 128 0 -1 396
box 8 4 76 44
use welltap_svt  __well_tap__6
timestamp 1667968642
transform 1 0 104 0 -1 388
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  add_afa_57_6
timestamp 1667968642
transform 1 0 328 0 -1 404
box 8 4 140 84
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_57_6_anx
timestamp 1667968642
transform 1 0 208 0 -1 396
box 8 4 36 60
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_57_6_al
timestamp 1667968642
transform 1 0 248 0 -1 396
box 8 4 76 48
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_55_6
timestamp 1668056734
transform 1 0 472 0 -1 396
box 2 -1 90 54
use _0_0std_0_0cells_0_0FAX1  add_afa_52_6
timestamp 1667968642
transform 1 0 560 0 -1 404
box 8 4 140 84
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_52_6_al
timestamp 1667968642
transform 1 0 712 0 -1 396
box 8 4 76 48
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_52_6
timestamp 1667968642
transform 1 0 856 0 -1 396
box 8 4 76 44
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_52_6
timestamp 1667968642
transform 1 0 792 0 -1 392
box 8 4 28 36
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_52_6
timestamp 1668054752
transform 1 0 824 0 -1 392
box 3 -1 28 37
use welltap_svt  __well_tap__7
timestamp 1667968642
transform 1 0 944 0 -1 388
box 8 4 12 24
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_57_6
timestamp 1667968642
transform 1 0 128 0 1 416
box 8 4 28 36
use welltap_svt  __well_tap__8
timestamp 1667968642
transform 1 0 104 0 1 420
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_57_6
timestamp 1668056734
transform 1 0 160 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0FAX1  add_afa_56_6
timestamp 1667968642
transform 1 0 336 0 1 404
box 8 4 140 84
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_57_6
timestamp 1668056734
transform 1 0 248 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_57_6
timestamp 1668056734
transform 1 0 480 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_52_6
timestamp 1668056734
transform 1 0 568 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_52_6
timestamp 1668056734
transform 1 0 656 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_52_6
timestamp 1668056734
transform 1 0 744 0 1 412
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_52_6
timestamp 1668056734
transform 1 0 832 0 1 412
box 2 -1 90 54
use welltap_svt  __well_tap__9
timestamp 1667968642
transform 1 0 944 0 1 420
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1667968642
transform 1 0 104 0 -1 564
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_57_6
timestamp 1668054752
transform 1 0 128 0 -1 568
box 3 -1 28 37
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_57_6
timestamp 1668056734
transform 1 0 160 0 -1 572
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_56_6
timestamp 1668056734
transform 1 0 336 0 -1 572
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_56_6
timestamp 1668056734
transform 1 0 248 0 -1 572
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_56_6_al
timestamp 1667968642
transform 1 0 432 0 -1 572
box 8 4 76 48
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_56_6_anx
timestamp 1667968642
transform 1 0 520 0 -1 572
box 8 4 36 60
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_51_6
timestamp 1668056734
transform 1 0 568 0 -1 572
box 2 -1 90 54
use _0_0std_0_0cells_0_0FAX1  add_afa_51_6
timestamp 1667968642
transform 1 0 664 0 -1 580
box 8 4 140 84
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_51_6_al
timestamp 1667968642
transform 1 0 816 0 -1 572
box 8 4 76 48
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_51_6_anx
timestamp 1667968642
transform 1 0 896 0 -1 572
box 8 4 36 60
use welltap_svt  __well_tap__11
timestamp 1667968642
transform 1 0 944 0 -1 564
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1667968642
transform 1 0 104 0 1 588
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_adel_adelay_52_6
timestamp 1668054752
transform 1 0 160 0 1 584
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_adel_adelay_51_6
timestamp 1668054752
transform 1 0 128 0 1 584
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_adel_adelay_50_6
timestamp 1668054752
transform 1 0 192 0 1 584
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_acinv
timestamp 1668054752
transform 1 0 224 0 1 584
box 3 -1 28 37
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_56_6
timestamp 1668056734
transform 1 0 256 0 1 580
box 2 -1 90 54
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_56_6
timestamp 1667968642
transform 1 0 464 0 1 584
box 8 4 28 36
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_56_6
timestamp 1668054752
transform 1 0 432 0 1 584
box 3 -1 28 37
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_56_6
timestamp 1668056734
transform 1 0 344 0 1 580
box 2 -1 90 54
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_56_6
timestamp 1667968642
transform 1 0 496 0 1 580
box 8 4 76 44
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_51_6
timestamp 1668056734
transform 1 0 576 0 1 580
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_51_6
timestamp 1668056734
transform 1 0 664 0 1 580
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  output_acopybuf_adatalatches_50_6
timestamp 1668056734
transform 1 0 664 0 -1 684
box 2 -1 90 54
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_51_6
timestamp 1667968642
transform 1 0 856 0 1 580
box 8 4 76 44
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_51_6
timestamp 1668056734
transform 1 0 760 0 1 580
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  ymerge_adatalatches_50_6
timestamp 1668056734
transform 1 0 752 0 -1 684
box 2 -1 90 54
use welltap_svt  __well_tap__13
timestamp 1667968642
transform 1 0 944 0 1 588
box 8 4 12 24
use _0_0std_0_0cells_0_0NAND2X1  ymerge_apg_apulsegen
timestamp 1667968642
transform 1 0 128 0 1 692
box 8 4 36 36
use _0_0std_0_0cells_0_0NOR2X1  ymerge_aoutgate
timestamp 1667968642
transform 1 0 200 0 1 696
box 8 4 36 40
use welltap_svt  __well_tap__14
timestamp 1667968642
transform 1 0 104 0 -1 676
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1667968642
transform 1 0 104 0 1 700
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_ainv1
timestamp 1668054752
transform 1 0 160 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_aoutgateinv
timestamp 1668054752
transform 1 0 168 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_ainv1
timestamp 1668054752
transform 1 0 128 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccB_adel_adelay_53_6
timestamp 1668054752
transform 1 0 192 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0NOR2X1  ymerge_amccB_aresetnor
timestamp 1667968642
transform 1 0 280 0 1 696
box 8 4 36 40
use _0_0std_0_0cells_0_0NOR2X1  ymerge_amccA_aresetnor
timestamp 1667968642
transform 1 0 320 0 1 696
box 8 4 36 40
use _0_0std_0_0cells_0_0NAND2X1  output_acopybuf_afcc_apg_apulsegen
timestamp 1667968642
transform 1 0 240 0 1 692
box 8 4 36 36
use _0_0std_0_0cells_0_0NOR2X1  yzero_acontrolgate
timestamp 1667968642
transform 1 0 224 0 -1 680
box 8 4 36 40
use _0_0cell_0_0gcelem3x0  ymerge_amccB_acelem_acx0
timestamp 1668055478
transform 1 0 264 0 -1 680
box 8 4 108 36
use _0_0std_0_0cells_0_0NAND2X1  ymerge_asplitB
timestamp 1667968642
transform 1 0 408 0 -1 684
box 8 4 36 36
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_acinv
timestamp 1668054752
transform 1 0 456 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_adel_adelay_52_6
timestamp 1668054752
transform 1 0 360 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_adel_adelay_51_6
timestamp 1668054752
transform 1 0 392 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_adel_adelay_50_6
timestamp 1668054752
transform 1 0 424 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_acB
timestamp 1668054752
transform 1 0 376 0 -1 680
box 3 -1 28 37
use _0_0cell_0_0gcelem3x0  ymerge_amccA_acelem_acx0
timestamp 1668055478
transform 1 0 448 0 -1 680
box 8 4 108 36
use _0_0std_0_0cells_0_0NAND2X1  ymerge_asplitA
timestamp 1667968642
transform 1 0 592 0 -1 684
box 8 4 36 36
use _0_0std_0_0cells_0_0NOR2X2  initialBuf_adatalatches_50_6_anx
timestamp 1667968642
transform 1 0 568 0 1 692
box 8 4 36 60
use _0_0std_0_0cells_0_0NOR2X1  initialBuf_afcc_aresetnor
timestamp 1667968642
transform 1 0 488 0 1 696
box 8 4 36 40
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_57_6
timestamp 1668054752
transform 1 0 528 0 1 696
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_acA
timestamp 1668054752
transform 1 0 560 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0FAX1  add_afa_50_6
timestamp 1667968642
transform 1 0 712 0 1 684
box 8 4 140 84
use _0_0std_0_0cells_0_0LATCHINV  initialBuf_adatalatches_50_6_al
timestamp 1667968642
transform 1 0 624 0 1 692
box 8 4 76 48
use _0_0std_0_0cells_0_0INVX1  ymerge_acbMaker
timestamp 1668054752
transform 1 0 632 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0MUX2X1  ymerge_amuxes_50_6
timestamp 1667968642
transform 1 0 856 0 1 692
box 8 4 76 44
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_50_6
timestamp 1668054752
transform 1 0 872 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amuxinv_51_6
timestamp 1668054752
transform 1 0 840 0 -1 680
box 3 -1 28 37
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_51_6
timestamp 1667968642
transform 1 0 904 0 -1 680
box 8 4 28 36
use welltap_svt  __well_tap__15
timestamp 1667968642
transform 1 0 944 0 -1 676
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1667968642
transform 1 0 944 0 1 700
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1667968642
transform 1 0 104 0 -1 816
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_adel_adelay_53_6
timestamp 1668054752
transform 1 0 192 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_adel_adelay_52_6
timestamp 1668054752
transform 1 0 160 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_adel_adelay_51_6
timestamp 1668054752
transform 1 0 128 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_ainv2
timestamp 1668054752
transform 1 0 256 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_adel_adelay_53_6
timestamp 1668054752
transform 1 0 288 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_adel_adelay_52_6
timestamp 1668054752
transform 1 0 320 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_ainv2
timestamp 1668054752
transform 1 0 224 0 -1 820
box 3 -1 28 37
use _0_0cell_0_0gcelem2x0  initialBuf_afcc_acelem_acx0
timestamp 1667972760
transform 1 0 416 0 -1 820
box 8 0 90 36
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_acinv
timestamp 1668054752
transform 1 0 384 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_amccA_adel_adelay_53_6
timestamp 1668054752
transform 1 0 352 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_56_6
timestamp 1668054752
transform 1 0 536 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_55_6
timestamp 1668054752
transform 1 0 568 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_54_6
timestamp 1668054752
transform 1 0 600 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_ainv1
timestamp 1668054752
transform 1 0 504 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesB_50_6
timestamp 1668056734
transform 1 0 720 0 -1 824
box 2 -1 90 54
use _0_0std_0_0cells_0_0LATCH  add_adatalatchesA_50_6
timestamp 1668056734
transform 1 0 632 0 -1 824
box 2 -1 90 54
use _0_0std_0_0cells_0_0TIELOX1  add_ainitialcarry
timestamp 1667968642
transform 1 0 864 0 -1 820
box 8 4 28 36
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_ainv1
timestamp 1668054752
transform 1 0 808 0 -1 820
box 3 -1 28 37
use _0_0std_0_0cells_0_0TIELOX1  yzero_atempt_50_6
timestamp 1667968642
transform 1 0 904 0 -1 820
box 8 4 28 36
use welltap_svt  __well_tap__19
timestamp 1667968642
transform 1 0 944 0 -1 816
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1667968642
transform 1 0 104 0 1 832
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  ymerge_apg_adel_adelay_50_6
timestamp 1668054752
transform 1 0 128 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_54_6
timestamp 1668054752
transform 1 0 192 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_53_6
timestamp 1668054752
transform 1 0 160 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_52_6
timestamp 1668054752
transform 1 0 128 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_51_6
timestamp 1668054752
transform 1 0 160 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_50_6
timestamp 1668054752
transform 1 0 192 0 1 828
box 3 -1 28 37
use _0_0cell_0_0gcelem2x0  add_ainputcelem_acelem_acx0
timestamp 1667972760
transform 1 0 288 0 -1 912
box 8 0 90 36
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_51_6
timestamp 1668054752
transform 1 0 256 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_50_6
timestamp 1668054752
transform 1 0 256 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_adel_adelay_51_6
timestamp 1668054752
transform 1 0 320 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_apg_adel_adelay_50_6
timestamp 1668054752
transform 1 0 288 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_56_6
timestamp 1668054752
transform 1 0 224 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_55_6
timestamp 1668054752
transform 1 0 224 0 -1 912
box 3 -1 28 37
use _0_0cell_0_0gcelem2x0  output_aacknowledgecelem_acelem_acx0
timestamp 1667972760
transform 1 0 440 0 -1 912
box 8 0 90 36
use _0_0cell_0_0gcelem2x0  output_acopybuf_afcc_acelem_acx0
timestamp 1667972760
transform 1 0 424 0 1 828
box 8 0 90 36
use _0_0std_0_0cells_0_0NOR2X1  output_acopybuf_afcc_aresetnor
timestamp 1667968642
transform 1 0 384 0 1 828
box 8 4 36 40
use _0_0std_0_0cells_0_0INVX1  add_ainputcelem_ainv
timestamp 1668054752
transform 1 0 376 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_aacknowledgecelem_ainv
timestamp 1668054752
transform 1 0 408 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  ymerge_adel_adelay_57_6
timestamp 1668054752
transform 1 0 352 0 1 828
box 3 -1 28 37
use _0_0cell_0_0gcelem2x0  add_afcc_acelem_acx0
timestamp 1667972760
transform 1 0 560 0 -1 912
box 8 0 90 36
use _0_0std_0_0cells_0_0NAND2X1  add_afcc_apg_apulsegen
timestamp 1667968642
transform 1 0 512 0 1 824
box 8 4 36 36
use _0_0std_0_0cells_0_0NOR2X1  add_afcc_aresetnor
timestamp 1667968642
transform 1 0 584 0 1 828
box 8 4 36 40
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_acinv
timestamp 1668054752
transform 1 0 552 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_acinv
timestamp 1668054752
transform 1 0 528 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_53_6
timestamp 1668054752
transform 1 0 624 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_52_6
timestamp 1668054752
transform 1 0 656 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_51_6
timestamp 1668054752
transform 1 0 688 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_adel_adelay_50_6
timestamp 1668054752
transform 1 0 712 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_adel_adelay_52_6
timestamp 1668054752
transform 1 0 720 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_ainv2
timestamp 1668054752
transform 1 0 648 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_adel_adelay_53_6
timestamp 1668054752
transform 1 0 680 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0NAND2X1  initialBuf_afcc_apg_apulsegen
timestamp 1667968642
transform 1 0 816 0 1 824
box 8 4 36 36
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_53_6
timestamp 1668054752
transform 1 0 872 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_ainv2
timestamp 1668054752
transform 1 0 784 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_adel_adelay_53_6
timestamp 1668054752
transform 1 0 752 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_adel_adelay_51_6
timestamp 1668054752
transform 1 0 744 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  initialBuf_afcc_apg_adel_adelay_50_6
timestamp 1668054752
transform 1 0 776 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_57_6
timestamp 1668054752
transform 1 0 856 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_55_6
timestamp 1668054752
transform 1 0 808 0 -1 912
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_54_6
timestamp 1668054752
transform 1 0 840 0 -1 912
box 3 -1 28 37
use welltap_svt  __well_tap__21
timestamp 1667968642
transform 1 0 944 0 1 832
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_56_6
timestamp 1668054752
transform 1 0 888 0 1 828
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_52_6
timestamp 1668054752
transform 1 0 904 0 -1 912
box 3 -1 28 37
use welltap_svt  __well_tap__22
timestamp 1667968642
transform 1 0 104 0 -1 908
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1667968642
transform 1 0 104 0 1 932
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_52_6
timestamp 1668054752
transform 1 0 208 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_55_6
timestamp 1668054752
transform 1 0 304 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_54_6
timestamp 1668054752
transform 1 0 272 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_53_6
timestamp 1668054752
transform 1 0 240 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_adel_adelay_50_6
timestamp 1668054752
transform 1 0 464 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_57_6
timestamp 1668054752
transform 1 0 408 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  output_acopybuf_afcc_adel_adelay_56_6
timestamp 1668054752
transform 1 0 352 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_adel_adelay_52_6
timestamp 1668054752
transform 1 0 592 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_apg_adel_adelay_51_6
timestamp 1668054752
transform 1 0 528 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_57_6
timestamp 1668054752
transform 1 0 720 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_56_6
timestamp 1668054752
transform 1 0 656 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_51_6
timestamp 1668054752
transform 1 0 856 0 1 928
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_adelay_adelay_50_6
timestamp 1668054752
transform 1 0 784 0 1 928
box 3 -1 28 37
use welltap_svt  __well_tap__23
timestamp 1667968642
transform 1 0 944 0 -1 908
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1667968642
transform 1 0 944 0 1 932
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  add_afcc_alainv
timestamp 1668054752
transform 1 0 904 0 1 928
box 3 -1 28 37
use welltap_svt  __well_tap__26
timestamp 1667968642
transform 1 0 104 0 -1 996
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_51_6
timestamp 1668054752
transform 1 0 584 0 -1 1000
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_50_6
timestamp 1668054752
transform 1 0 536 0 -1 1000
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_53_6
timestamp 1668054752
transform 1 0 688 0 -1 1000
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_52_6
timestamp 1668054752
transform 1 0 632 0 -1 1000
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_55_6
timestamp 1668054752
transform 1 0 800 0 -1 1000
box 3 -1 28 37
use _0_0std_0_0cells_0_0INVX1  add_afcc_adel_adelay_54_6
timestamp 1668054752
transform 1 0 744 0 -1 1000
box 3 -1 28 37
use welltap_svt  __well_tap__27
timestamp 1667968642
transform 1 0 944 0 -1 996
box 8 4 12 24
<< labels >>
rlabel m2 s 982 920 984 928 6 L.d[0]
port 0 nsew signal input
rlabel m2 s 982 748 984 756 6 L.d[1]
port 1 nsew signal input
rlabel m2 s 982 492 984 500 6 L.d[2]
port 2 nsew signal input
rlabel m2 s 982 240 984 248 6 L.d[3]
port 3 nsew signal input
rlabel m2 s 80 304 82 312 6 L.d[4]
port 4 nsew signal input
rlabel m2 s 80 380 82 388 6 L.d[5]
port 5 nsew signal input
rlabel m2 s 80 616 82 624 6 L.d[6]
port 6 nsew signal input
rlabel m2 s 80 536 82 544 6 L.d[7]
port 7 nsew signal input
rlabel m2 s 80 928 82 936 6 L.r
port 8 nsew signal input
rlabel m2 s 756 1006 764 1008 6 L.a
port 9 nsew signal tristate
rlabel m2 s 982 324 984 332 6 C.d[0]
port 10 nsew signal input
rlabel m2 s 80 772 82 780 6 C.r
port 11 nsew signal input
rlabel m2 s 80 848 82 856 6 C.a
port 12 nsew signal tristate
rlabel m2 s 982 832 984 840 6 R.d[0]
port 13 nsew signal tristate
rlabel m2 s 982 664 984 672 6 R.d[1]
port 14 nsew signal tristate
rlabel m2 s 982 408 984 416 6 R.d[2]
port 15 nsew signal tristate
rlabel m2 s 982 152 984 160 6 R.d[3]
port 16 nsew signal tristate
rlabel m2 s 80 148 82 156 6 R.d[4]
port 17 nsew signal tristate
rlabel m2 s 80 224 82 232 6 R.d[5]
port 18 nsew signal tristate
rlabel m2 s 80 692 82 700 6 R.d[6]
port 19 nsew signal tristate
rlabel m2 s 80 460 82 468 6 R.d[7]
port 20 nsew signal tristate
rlabel m2 s 300 1006 308 1008 6 R.r
port 21 nsew signal tristate
rlabel m2 s 532 1006 540 1008 6 R.a
port 22 nsew signal input
rlabel m2 s 982 580 984 588 6 Reset
port 23 nsew signal input
<< end >>
