magic
tech sky130l
timestamp 1667968642
<< m1 >>
rect 8 80 12 84
rect 40 80 44 84
rect 72 80 76 84
rect 104 80 108 84
rect 136 80 140 84
rect 8 24 135 63
rect 8 4 12 8
rect 72 4 76 8
<< labels >>
rlabel m1 s 8 80 12 84 6 A
port 1 nsew signal input
rlabel m1 s 40 80 44 84 6 B
port 2 nsew signal input
rlabel m1 s 72 80 76 84 6 C
port 3 nsew signal input
rlabel m1 s 8 4 12 8 6 YC
port 4 nsew signal output
rlabel m1 s 72 4 76 8 6 YS
port 5 nsew signal output
rlabel m1 s 104 80 108 84 6 Vdd
port 6 nsew power input
rlabel m1 s 136 80 140 84 6 GND
port 7 nsew ground input
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 144 88
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
